-- Copyright (C) 1991-2009 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 9.0 Build 235 06/17/2009 Service Pack 2 SJ Web Edition
-- Created on Fri May 26 22:19:53 2017

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY UFC IS
    PORT (
        clock : IN STD_LOGIC;
        I : IN STD_LOGIC := '0';
        C : IN STD_LOGIC := '0';
        LD : OUT STD_LOGIC;
        CLS : OUT STD_LOGIC
    );
END UFC;

ARCHITECTURE BEHAVIOR OF UFC IS
    TYPE type_fstate IS (zero,one,two,three_CLS,four,five,seven_LD_CLS,eight,nine,fifteen_CLS);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,I,C)
    BEGIN
		LD <= '0';
		CLS <= '0';
		CASE fstate IS
			WHEN zero =>
				IF ((I = '1')) THEN
					reg_fstate <= one;
				ELSIF ((NOT((I = '1')) AND (C = '1'))) THEN
					reg_fstate <= fifteen_CLS;
				-- Inserting 'else' block to prevent latch inference
				ELSE
					reg_fstate <= zero;
				END IF;
			WHEN one =>
				IF (NOT((I = '1'))) THEN
					reg_fstate <= two;
				-- Inserting 'else' block to prevent latch inference
				ELSE
					reg_fstate <= one;
				END IF;
			WHEN two =>
				IF (((I = '1') AND NOT((C = '1')))) THEN
					reg_fstate <= three_CLS;
				ELSIF ((C = '1')) THEN
					reg_fstate <= fifteen_CLS;
				-- Inserting 'else' block to prevent latch inference
				ELSE
					reg_fstate <= two;
				END IF;
			WHEN three_CLS =>
				reg_fstate <= four;

				CLS <= '1';
			WHEN four =>
				IF (NOT((I = '1'))) THEN
					reg_fstate <= five;
				-- Inserting 'else' block to prevent latch inference
				ELSE
					reg_fstate <= four;
				END IF;
			WHEN five =>
				IF (((I = '1') AND NOT((C = '1')))) THEN
					reg_fstate <= seven_LD_CLS;
				ELSIF ((C = '1')) THEN
					reg_fstate <= fifteen_CLS;
				-- Inserting 'else' block to prevent latch inference
				ELSE
					reg_fstate <= five;
				END IF;
			WHEN seven_LD_CLS =>
				reg_fstate <= eight;

				CLS <= '1';

				LD <= '1';
			WHEN eight =>
				IF (NOT((I = '1'))) THEN
					reg_fstate <= nine;
				-- Inserting 'else' block to prevent latch inference
				ELSE
					reg_fstate <= eight;
				END IF;
			WHEN nine =>
				IF ((I = '1')) THEN
					reg_fstate <= seven_LD_CLS;
				ELSIF ((NOT((I = '1')) AND (C = '1'))) THEN
					reg_fstate <= fifteen_CLS;
				-- Inserting 'else' block to prevent latch inference
				ELSE
					reg_fstate <= nine;
				END IF;
			WHEN fifteen_CLS =>
				reg_fstate <= zero;

				CLS <= '1';
			WHEN OTHERS => 
				LD <= 'X';
				CLS <= 'X';
				report "Reach undefined state";
		END CASE;
    END PROCESS;
END BEHAVIOR;
