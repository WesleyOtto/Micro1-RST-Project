-- Copyright (C) 1991-2009 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 9.0 Build 235 06/17/2009 Service Pack 2 SJ Web Edition
-- Created on Fri May 20 21:49:41 2016

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY compfase2 IS
    PORT (
        CL : IN STD_LOGIC := '0';
        CK : IN STD_LOGIC;
        RealFase1 : OUT STD_LOGIC;
        RealFase2 : OUT STD_LOGIC
    );
END compfase2;

ARCHITECTURE BEHAVIOR OF compfase2 IS
    TYPE type_fstate IS (state1,state2,state3);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (CK,CL,reg_fstate)
    BEGIN
        IF (CL='1') THEN
            fstate <= state1;
        ELSIF (CK='1' AND CK'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate)
    BEGIN
        RealFase1 <= '0';
        RealFase2 <= '0';
        CASE fstate IS
            WHEN state1 =>
                reg_fstate <= state2;

                RealFase2 <= '0';

                RealFase1 <= '0';
            WHEN state2 =>
                reg_fstate <= state3;

                RealFase2 <= '1';

                RealFase1 <= '0';
            WHEN state3 =>
                reg_fstate <= state1;

                RealFase2 <= '0';

                RealFase1 <= '1';
            WHEN OTHERS => 
                RealFase1 <= 'X';
                RealFase2 <= 'X';
                report "Reach undefined state";
        END CASE;
    END PROCESS;
END BEHAVIOR;
