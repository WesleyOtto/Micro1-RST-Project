-- Copyright (C) 1991-2009 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 9.0 Build 235 06/17/2009 Service Pack 2 SJ Web Edition
-- Created on Fri May 13 23:58:10 2016

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY compfase IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        output1 : OUT STD_LOGIC;
        output2 : OUT STD_LOGIC
    );
END compfase;

ARCHITECTURE BEHAVIOR OF compfase IS
    TYPE type_fstate IS (state1,state2,state3,state4,state5,state6);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reset,reg_fstate)
    BEGIN
        IF (reset='1') THEN
            fstate <= state1;
        ELSIF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate)
    BEGIN
        output1 <= '0';
        output2 <= '0';
        CASE fstate IS
            WHEN state1 =>
                reg_fstate <= state2;
            WHEN state2 =>
                reg_fstate <= state3;

                output2 <= '1';
            WHEN state3 =>
                reg_fstate <= state4;

                output2 <= '1';
            WHEN state4 =>
                reg_fstate <= state5;

                output1 <= '1';
            WHEN state5 =>
                reg_fstate <= state6;

                output1 <= '1';
            WHEN state6 =>
                reg_fstate <= state1;
            WHEN OTHERS => 
                output1 <= 'X';
                output2 <= 'X';
                report "Reach undefined state";
        END CASE;
    END PROCESS;
END BEHAVIOR;
