-- Copyright (C) 1991-2009 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 9.0 Build 235 06/17/2009 Service Pack 2 SJ Web Edition
-- Created on Fri May 06 22:17:22 2016

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY UCF IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        E : IN STD_LOGIC := '0';
        C : IN STD_LOGIC := '0';
        Ld : OUT STD_LOGIC;
        Cls : OUT STD_LOGIC
    );
END UCF;

ARCHITECTURE BEHAVIOR OF UCF IS
    TYPE type_fstate IS (Zero,Um,Dois,Tres,Quatro,Cinco,Sete_LD_CL,Oito,Nove,Quinze);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,E,C)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= Zero;
            Ld <= '0';
            Cls <= '0';
        ELSE
            Ld <= '0';
            Cls <= '0';
            CASE fstate IS
                WHEN Zero =>
                    IF ((E = '1')) THEN
                        reg_fstate <= Um;
                    ELSIF ((NOT((E = '1')) AND (C = '1'))) THEN
                        reg_fstate <= Quinze;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Zero;
                    END IF;
                WHEN Um =>
                    IF (NOT((E = '1'))) THEN
                        reg_fstate <= Dois;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Um;
                    END IF;
                WHEN Dois =>
                    IF ((E = '1')) THEN
                        reg_fstate <= Tres;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Dois;
                    END IF;
                WHEN Tres =>
                    reg_fstate <= Quatro;

                    Cls <= '1';
                WHEN Quatro =>
                    IF (NOT((E = '1'))) THEN
                        reg_fstate <= Cinco;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Quatro;
                    END IF;
                WHEN Cinco =>
                    IF ((E = '1')) THEN
                        reg_fstate <= Sete_LD_CL;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Cinco;
                    END IF;
                WHEN Sete_LD_CL =>
                    reg_fstate <= Oito;

                    Ld <= '1';

                    Cls <= '1';
                WHEN Oito =>
                    IF (NOT((E = '1'))) THEN
                        reg_fstate <= Nove;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Oito;
                    END IF;
                WHEN Nove =>
                    IF ((E = '1')) THEN
                        reg_fstate <= Sete_LD_CL;
                    ELSIF ((NOT((E = '1')) AND (C = '1'))) THEN
                        reg_fstate <= Quinze;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Nove;
                    END IF;
                WHEN Quinze =>
                    reg_fstate <= Zero;

                    Cls <= '1';
                WHEN OTHERS => 
                    Ld <= 'X';
                    Cls <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
